` include "adder_subtractor"
module bcd_adder(
    input [0:3] a,b,
    output [0:3] sum
)