module hellow();
initial begin
	$display("hellow world");
end
endmodule
